
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h76713fc1;
    ram_cell[       1] = 32'h0;  // 32'hb41015fe;
    ram_cell[       2] = 32'h0;  // 32'hca69b7fb;
    ram_cell[       3] = 32'h0;  // 32'h4815070d;
    ram_cell[       4] = 32'h0;  // 32'h0db5b39f;
    ram_cell[       5] = 32'h0;  // 32'h26075227;
    ram_cell[       6] = 32'h0;  // 32'h197b362d;
    ram_cell[       7] = 32'h0;  // 32'h125214ff;
    ram_cell[       8] = 32'h0;  // 32'hd0bef1c2;
    ram_cell[       9] = 32'h0;  // 32'h3844a5c2;
    ram_cell[      10] = 32'h0;  // 32'h7448c059;
    ram_cell[      11] = 32'h0;  // 32'hf9338dee;
    ram_cell[      12] = 32'h0;  // 32'h3e948e9d;
    ram_cell[      13] = 32'h0;  // 32'hd96df32f;
    ram_cell[      14] = 32'h0;  // 32'h375a584c;
    ram_cell[      15] = 32'h0;  // 32'h1766c95c;
    ram_cell[      16] = 32'h0;  // 32'h4b866acf;
    ram_cell[      17] = 32'h0;  // 32'h9e431577;
    ram_cell[      18] = 32'h0;  // 32'h717c9a21;
    ram_cell[      19] = 32'h0;  // 32'h48f2f9e4;
    ram_cell[      20] = 32'h0;  // 32'heaa2dc0a;
    ram_cell[      21] = 32'h0;  // 32'hb568e8bd;
    ram_cell[      22] = 32'h0;  // 32'h8a01f686;
    ram_cell[      23] = 32'h0;  // 32'h91c719ad;
    ram_cell[      24] = 32'h0;  // 32'hc2a02371;
    ram_cell[      25] = 32'h0;  // 32'h75557758;
    ram_cell[      26] = 32'h0;  // 32'h7e242138;
    ram_cell[      27] = 32'h0;  // 32'h0d4f5d79;
    ram_cell[      28] = 32'h0;  // 32'hb3872a15;
    ram_cell[      29] = 32'h0;  // 32'hadbed708;
    ram_cell[      30] = 32'h0;  // 32'hb12013bd;
    ram_cell[      31] = 32'h0;  // 32'h514cbd18;
    ram_cell[      32] = 32'h0;  // 32'h568e4051;
    ram_cell[      33] = 32'h0;  // 32'h9815294e;
    ram_cell[      34] = 32'h0;  // 32'h2dbb00e8;
    ram_cell[      35] = 32'h0;  // 32'h16c30ec3;
    ram_cell[      36] = 32'h0;  // 32'h651ba4de;
    ram_cell[      37] = 32'h0;  // 32'h10777bcd;
    ram_cell[      38] = 32'h0;  // 32'hcd790f0e;
    ram_cell[      39] = 32'h0;  // 32'h0765c601;
    ram_cell[      40] = 32'h0;  // 32'h09133fd7;
    ram_cell[      41] = 32'h0;  // 32'hcef91ef7;
    ram_cell[      42] = 32'h0;  // 32'hdc60d457;
    ram_cell[      43] = 32'h0;  // 32'h0ea64981;
    ram_cell[      44] = 32'h0;  // 32'he012daba;
    ram_cell[      45] = 32'h0;  // 32'h1dd75389;
    ram_cell[      46] = 32'h0;  // 32'h7c56966b;
    ram_cell[      47] = 32'h0;  // 32'he9019f25;
    ram_cell[      48] = 32'h0;  // 32'h315bb35c;
    ram_cell[      49] = 32'h0;  // 32'h37a14294;
    ram_cell[      50] = 32'h0;  // 32'hf38015d6;
    ram_cell[      51] = 32'h0;  // 32'hd27567e8;
    ram_cell[      52] = 32'h0;  // 32'h7353335c;
    ram_cell[      53] = 32'h0;  // 32'hd8a9cd9b;
    ram_cell[      54] = 32'h0;  // 32'h0ee4dea4;
    ram_cell[      55] = 32'h0;  // 32'h56bbf621;
    ram_cell[      56] = 32'h0;  // 32'hd6d69e53;
    ram_cell[      57] = 32'h0;  // 32'hfe8f81fa;
    ram_cell[      58] = 32'h0;  // 32'hb2712993;
    ram_cell[      59] = 32'h0;  // 32'h33020894;
    ram_cell[      60] = 32'h0;  // 32'h6fecf6a0;
    ram_cell[      61] = 32'h0;  // 32'he0496dda;
    ram_cell[      62] = 32'h0;  // 32'h7ac55f44;
    ram_cell[      63] = 32'h0;  // 32'h882213f2;
    ram_cell[      64] = 32'h0;  // 32'hd34ae3bb;
    ram_cell[      65] = 32'h0;  // 32'hab3da0fb;
    ram_cell[      66] = 32'h0;  // 32'h6835aa2b;
    ram_cell[      67] = 32'h0;  // 32'h2f6d0d78;
    ram_cell[      68] = 32'h0;  // 32'h7cd0d18b;
    ram_cell[      69] = 32'h0;  // 32'he227882e;
    ram_cell[      70] = 32'h0;  // 32'hda88fd29;
    ram_cell[      71] = 32'h0;  // 32'hb9a86ea8;
    ram_cell[      72] = 32'h0;  // 32'hba087f8d;
    ram_cell[      73] = 32'h0;  // 32'h0c6a2e7e;
    ram_cell[      74] = 32'h0;  // 32'hc67638c8;
    ram_cell[      75] = 32'h0;  // 32'hfb0e8d27;
    ram_cell[      76] = 32'h0;  // 32'h3508cf6e;
    ram_cell[      77] = 32'h0;  // 32'hf52cff64;
    ram_cell[      78] = 32'h0;  // 32'h123b5ab7;
    ram_cell[      79] = 32'h0;  // 32'he9742fa7;
    ram_cell[      80] = 32'h0;  // 32'h5aac6d6e;
    ram_cell[      81] = 32'h0;  // 32'he228a949;
    ram_cell[      82] = 32'h0;  // 32'h6cc0190c;
    ram_cell[      83] = 32'h0;  // 32'he1739c7d;
    ram_cell[      84] = 32'h0;  // 32'had377249;
    ram_cell[      85] = 32'h0;  // 32'ha36b7e39;
    ram_cell[      86] = 32'h0;  // 32'h5c53b475;
    ram_cell[      87] = 32'h0;  // 32'h7408d3e3;
    ram_cell[      88] = 32'h0;  // 32'h209522a3;
    ram_cell[      89] = 32'h0;  // 32'h95e6c98b;
    ram_cell[      90] = 32'h0;  // 32'haaab7085;
    ram_cell[      91] = 32'h0;  // 32'h22f83e36;
    ram_cell[      92] = 32'h0;  // 32'he7e3850a;
    ram_cell[      93] = 32'h0;  // 32'ha41ea60a;
    ram_cell[      94] = 32'h0;  // 32'hb744e0a9;
    ram_cell[      95] = 32'h0;  // 32'hfb7ae13f;
    ram_cell[      96] = 32'h0;  // 32'hc770d8e4;
    ram_cell[      97] = 32'h0;  // 32'h970b6f30;
    ram_cell[      98] = 32'h0;  // 32'h923f8b71;
    ram_cell[      99] = 32'h0;  // 32'hfe3df851;
    ram_cell[     100] = 32'h0;  // 32'hf697abcd;
    ram_cell[     101] = 32'h0;  // 32'haa302934;
    ram_cell[     102] = 32'h0;  // 32'hd473d3bf;
    ram_cell[     103] = 32'h0;  // 32'h4b341ce5;
    ram_cell[     104] = 32'h0;  // 32'hf5e68a1e;
    ram_cell[     105] = 32'h0;  // 32'h14a1cbe5;
    ram_cell[     106] = 32'h0;  // 32'hbe43870b;
    ram_cell[     107] = 32'h0;  // 32'h1e3ff3b0;
    ram_cell[     108] = 32'h0;  // 32'h5ec52bdf;
    ram_cell[     109] = 32'h0;  // 32'h0b50ce91;
    ram_cell[     110] = 32'h0;  // 32'hea015cc7;
    ram_cell[     111] = 32'h0;  // 32'hb4592198;
    ram_cell[     112] = 32'h0;  // 32'h9b027d71;
    ram_cell[     113] = 32'h0;  // 32'h6fe1278f;
    ram_cell[     114] = 32'h0;  // 32'h1ae0c279;
    ram_cell[     115] = 32'h0;  // 32'h22bfb706;
    ram_cell[     116] = 32'h0;  // 32'hb61335a8;
    ram_cell[     117] = 32'h0;  // 32'haf627d50;
    ram_cell[     118] = 32'h0;  // 32'hf12f5994;
    ram_cell[     119] = 32'h0;  // 32'he1dfb453;
    ram_cell[     120] = 32'h0;  // 32'h13b89e65;
    ram_cell[     121] = 32'h0;  // 32'ha1a27645;
    ram_cell[     122] = 32'h0;  // 32'hf2a1fcb8;
    ram_cell[     123] = 32'h0;  // 32'h913984c6;
    ram_cell[     124] = 32'h0;  // 32'h9ce29da5;
    ram_cell[     125] = 32'h0;  // 32'hf0490a95;
    ram_cell[     126] = 32'h0;  // 32'hd0113e96;
    ram_cell[     127] = 32'h0;  // 32'h901e12a3;
    ram_cell[     128] = 32'h0;  // 32'h76eb5b0d;
    ram_cell[     129] = 32'h0;  // 32'h9ecf9e06;
    ram_cell[     130] = 32'h0;  // 32'hc3112965;
    ram_cell[     131] = 32'h0;  // 32'h7b99c46e;
    ram_cell[     132] = 32'h0;  // 32'he01b6384;
    ram_cell[     133] = 32'h0;  // 32'h2cf1bda7;
    ram_cell[     134] = 32'h0;  // 32'h7722b33c;
    ram_cell[     135] = 32'h0;  // 32'h8f087b29;
    ram_cell[     136] = 32'h0;  // 32'ha82b7538;
    ram_cell[     137] = 32'h0;  // 32'h7fe64f01;
    ram_cell[     138] = 32'h0;  // 32'h36cbe5a7;
    ram_cell[     139] = 32'h0;  // 32'ha7f96baa;
    ram_cell[     140] = 32'h0;  // 32'hfaeca288;
    ram_cell[     141] = 32'h0;  // 32'h2328b9c2;
    ram_cell[     142] = 32'h0;  // 32'hc5b714eb;
    ram_cell[     143] = 32'h0;  // 32'h5299152e;
    ram_cell[     144] = 32'h0;  // 32'h0a9ac926;
    ram_cell[     145] = 32'h0;  // 32'he4b9b010;
    ram_cell[     146] = 32'h0;  // 32'h78793348;
    ram_cell[     147] = 32'h0;  // 32'hfa921e09;
    ram_cell[     148] = 32'h0;  // 32'hc6cf413c;
    ram_cell[     149] = 32'h0;  // 32'he8cdd3dd;
    ram_cell[     150] = 32'h0;  // 32'hf6364d5a;
    ram_cell[     151] = 32'h0;  // 32'heaaf637b;
    ram_cell[     152] = 32'h0;  // 32'hf070e95c;
    ram_cell[     153] = 32'h0;  // 32'hd9e048c0;
    ram_cell[     154] = 32'h0;  // 32'h40553cba;
    ram_cell[     155] = 32'h0;  // 32'h3fff6286;
    ram_cell[     156] = 32'h0;  // 32'ha2e20f14;
    ram_cell[     157] = 32'h0;  // 32'h7bd564dd;
    ram_cell[     158] = 32'h0;  // 32'h571f5d55;
    ram_cell[     159] = 32'h0;  // 32'h9e954a7a;
    ram_cell[     160] = 32'h0;  // 32'h54f11b53;
    ram_cell[     161] = 32'h0;  // 32'hf2b2f306;
    ram_cell[     162] = 32'h0;  // 32'h070df207;
    ram_cell[     163] = 32'h0;  // 32'he41cf727;
    ram_cell[     164] = 32'h0;  // 32'h722c55fd;
    ram_cell[     165] = 32'h0;  // 32'hec19e20e;
    ram_cell[     166] = 32'h0;  // 32'hf31fa61e;
    ram_cell[     167] = 32'h0;  // 32'h837e0bd0;
    ram_cell[     168] = 32'h0;  // 32'hc72ed7cd;
    ram_cell[     169] = 32'h0;  // 32'h64ca28f2;
    ram_cell[     170] = 32'h0;  // 32'hc58c7f4e;
    ram_cell[     171] = 32'h0;  // 32'hd18b780d;
    ram_cell[     172] = 32'h0;  // 32'he58ea5d6;
    ram_cell[     173] = 32'h0;  // 32'hbd713a22;
    ram_cell[     174] = 32'h0;  // 32'hd0b190eb;
    ram_cell[     175] = 32'h0;  // 32'he562b050;
    ram_cell[     176] = 32'h0;  // 32'hcb2d7a9e;
    ram_cell[     177] = 32'h0;  // 32'h8cecc288;
    ram_cell[     178] = 32'h0;  // 32'hc1a57e45;
    ram_cell[     179] = 32'h0;  // 32'h09156ef2;
    ram_cell[     180] = 32'h0;  // 32'h768f7da9;
    ram_cell[     181] = 32'h0;  // 32'h702f68f3;
    ram_cell[     182] = 32'h0;  // 32'h87369437;
    ram_cell[     183] = 32'h0;  // 32'hf20e9aea;
    ram_cell[     184] = 32'h0;  // 32'h4143481e;
    ram_cell[     185] = 32'h0;  // 32'h0b3773d0;
    ram_cell[     186] = 32'h0;  // 32'h70c09188;
    ram_cell[     187] = 32'h0;  // 32'h56ce9a52;
    ram_cell[     188] = 32'h0;  // 32'hd67b3ad7;
    ram_cell[     189] = 32'h0;  // 32'ha66e816d;
    ram_cell[     190] = 32'h0;  // 32'ha39a070a;
    ram_cell[     191] = 32'h0;  // 32'h5804230c;
    ram_cell[     192] = 32'h0;  // 32'hfd90a837;
    ram_cell[     193] = 32'h0;  // 32'h3482d074;
    ram_cell[     194] = 32'h0;  // 32'h155338e9;
    ram_cell[     195] = 32'h0;  // 32'h4847adcf;
    ram_cell[     196] = 32'h0;  // 32'h3d43fefd;
    ram_cell[     197] = 32'h0;  // 32'h8a5285b1;
    ram_cell[     198] = 32'h0;  // 32'h758202cf;
    ram_cell[     199] = 32'h0;  // 32'h8680c635;
    ram_cell[     200] = 32'h0;  // 32'hf5e32cef;
    ram_cell[     201] = 32'h0;  // 32'he42125b1;
    ram_cell[     202] = 32'h0;  // 32'hec08e67f;
    ram_cell[     203] = 32'h0;  // 32'h0a83edf5;
    ram_cell[     204] = 32'h0;  // 32'h42c3e498;
    ram_cell[     205] = 32'h0;  // 32'h51b7ee15;
    ram_cell[     206] = 32'h0;  // 32'h077c8dbd;
    ram_cell[     207] = 32'h0;  // 32'ha231f998;
    ram_cell[     208] = 32'h0;  // 32'h944fef38;
    ram_cell[     209] = 32'h0;  // 32'h2d064355;
    ram_cell[     210] = 32'h0;  // 32'ha88b0910;
    ram_cell[     211] = 32'h0;  // 32'h63f2c540;
    ram_cell[     212] = 32'h0;  // 32'h9f201a3f;
    ram_cell[     213] = 32'h0;  // 32'h64efd340;
    ram_cell[     214] = 32'h0;  // 32'hda790d5a;
    ram_cell[     215] = 32'h0;  // 32'h3b5a63cc;
    ram_cell[     216] = 32'h0;  // 32'h856f0588;
    ram_cell[     217] = 32'h0;  // 32'h33df090c;
    ram_cell[     218] = 32'h0;  // 32'h2983c1c7;
    ram_cell[     219] = 32'h0;  // 32'h62d161bd;
    ram_cell[     220] = 32'h0;  // 32'h1b2700b6;
    ram_cell[     221] = 32'h0;  // 32'h4434debe;
    ram_cell[     222] = 32'h0;  // 32'he4948649;
    ram_cell[     223] = 32'h0;  // 32'h36dec246;
    ram_cell[     224] = 32'h0;  // 32'h7295cccd;
    ram_cell[     225] = 32'h0;  // 32'hb0b4b0ea;
    ram_cell[     226] = 32'h0;  // 32'h932dfc0f;
    ram_cell[     227] = 32'h0;  // 32'h90c9c4d4;
    ram_cell[     228] = 32'h0;  // 32'hf0c0724d;
    ram_cell[     229] = 32'h0;  // 32'h48686cf3;
    ram_cell[     230] = 32'h0;  // 32'h32c53311;
    ram_cell[     231] = 32'h0;  // 32'hdcc5142f;
    ram_cell[     232] = 32'h0;  // 32'h7b44c677;
    ram_cell[     233] = 32'h0;  // 32'haeeb3bfc;
    ram_cell[     234] = 32'h0;  // 32'h9acbd2c7;
    ram_cell[     235] = 32'h0;  // 32'hbcd43b27;
    ram_cell[     236] = 32'h0;  // 32'h37c3b605;
    ram_cell[     237] = 32'h0;  // 32'h35f4aa7d;
    ram_cell[     238] = 32'h0;  // 32'h4497f459;
    ram_cell[     239] = 32'h0;  // 32'h47018c74;
    ram_cell[     240] = 32'h0;  // 32'he3bf8658;
    ram_cell[     241] = 32'h0;  // 32'hae07a5bb;
    ram_cell[     242] = 32'h0;  // 32'h87486145;
    ram_cell[     243] = 32'h0;  // 32'h264e8451;
    ram_cell[     244] = 32'h0;  // 32'hd2b18d32;
    ram_cell[     245] = 32'h0;  // 32'h1664faae;
    ram_cell[     246] = 32'h0;  // 32'hba08fa13;
    ram_cell[     247] = 32'h0;  // 32'hafe129b7;
    ram_cell[     248] = 32'h0;  // 32'h1acaace2;
    ram_cell[     249] = 32'h0;  // 32'ha1d325b5;
    ram_cell[     250] = 32'h0;  // 32'hc5993846;
    ram_cell[     251] = 32'h0;  // 32'h4be0730a;
    ram_cell[     252] = 32'h0;  // 32'h572e1900;
    ram_cell[     253] = 32'h0;  // 32'he798810f;
    ram_cell[     254] = 32'h0;  // 32'h6d9c3572;
    ram_cell[     255] = 32'h0;  // 32'h3af75cfd;
    // src matrix A
    ram_cell[     256] = 32'h4879ebee;
    ram_cell[     257] = 32'hbab3caba;
    ram_cell[     258] = 32'hc51c4a06;
    ram_cell[     259] = 32'hce1ab7de;
    ram_cell[     260] = 32'h54d88228;
    ram_cell[     261] = 32'ha6b50014;
    ram_cell[     262] = 32'h87778383;
    ram_cell[     263] = 32'h4860a4a9;
    ram_cell[     264] = 32'h09a54aa6;
    ram_cell[     265] = 32'h32ed8f56;
    ram_cell[     266] = 32'h949af197;
    ram_cell[     267] = 32'h8c18df5b;
    ram_cell[     268] = 32'h40603b4e;
    ram_cell[     269] = 32'ha685e0df;
    ram_cell[     270] = 32'h1f742e39;
    ram_cell[     271] = 32'hf71bbea6;
    ram_cell[     272] = 32'hb97d08ec;
    ram_cell[     273] = 32'hcf1a46e0;
    ram_cell[     274] = 32'h8db4b06e;
    ram_cell[     275] = 32'h48f6e7fd;
    ram_cell[     276] = 32'ha718e618;
    ram_cell[     277] = 32'h4df815c7;
    ram_cell[     278] = 32'h59b11a91;
    ram_cell[     279] = 32'ha1da327c;
    ram_cell[     280] = 32'h17442f15;
    ram_cell[     281] = 32'h77d2634e;
    ram_cell[     282] = 32'h0e1ff72e;
    ram_cell[     283] = 32'hfeed16e8;
    ram_cell[     284] = 32'hdd8b3ccc;
    ram_cell[     285] = 32'hf88de47a;
    ram_cell[     286] = 32'hd57e34f6;
    ram_cell[     287] = 32'h30019b15;
    ram_cell[     288] = 32'h7484d92f;
    ram_cell[     289] = 32'he29e59ad;
    ram_cell[     290] = 32'h1b5bdd07;
    ram_cell[     291] = 32'h37a15636;
    ram_cell[     292] = 32'h9e169e92;
    ram_cell[     293] = 32'hc372a972;
    ram_cell[     294] = 32'hc384e290;
    ram_cell[     295] = 32'ha0bb646b;
    ram_cell[     296] = 32'h99f25484;
    ram_cell[     297] = 32'h319bd4c6;
    ram_cell[     298] = 32'ha77a279e;
    ram_cell[     299] = 32'hc8ee436d;
    ram_cell[     300] = 32'h861956e0;
    ram_cell[     301] = 32'h942aee52;
    ram_cell[     302] = 32'hdb480828;
    ram_cell[     303] = 32'h3aec04f7;
    ram_cell[     304] = 32'h6705f29b;
    ram_cell[     305] = 32'heaa8824e;
    ram_cell[     306] = 32'hd529a8bf;
    ram_cell[     307] = 32'h6dd37dbb;
    ram_cell[     308] = 32'hd1c8349c;
    ram_cell[     309] = 32'h4ff8b174;
    ram_cell[     310] = 32'h1a0e2905;
    ram_cell[     311] = 32'he1477ca9;
    ram_cell[     312] = 32'hd154facc;
    ram_cell[     313] = 32'hf1bf357c;
    ram_cell[     314] = 32'h12858c5b;
    ram_cell[     315] = 32'ha6c3a2c9;
    ram_cell[     316] = 32'hf33cd0cd;
    ram_cell[     317] = 32'he47648f3;
    ram_cell[     318] = 32'h8a2e2ce7;
    ram_cell[     319] = 32'h16673371;
    ram_cell[     320] = 32'hc9403920;
    ram_cell[     321] = 32'h7031a2a0;
    ram_cell[     322] = 32'h6321b250;
    ram_cell[     323] = 32'h46c541b0;
    ram_cell[     324] = 32'h4b01ad4f;
    ram_cell[     325] = 32'hc286a943;
    ram_cell[     326] = 32'hc718605b;
    ram_cell[     327] = 32'hdd17fa36;
    ram_cell[     328] = 32'h832c377b;
    ram_cell[     329] = 32'h8d61f042;
    ram_cell[     330] = 32'h70679e6c;
    ram_cell[     331] = 32'h30c72604;
    ram_cell[     332] = 32'hbe4e677f;
    ram_cell[     333] = 32'hde4c13e2;
    ram_cell[     334] = 32'h69b35d43;
    ram_cell[     335] = 32'h04c234b1;
    ram_cell[     336] = 32'h852c5910;
    ram_cell[     337] = 32'h9b523ccc;
    ram_cell[     338] = 32'h050bd407;
    ram_cell[     339] = 32'h0003e8d4;
    ram_cell[     340] = 32'hd15d748a;
    ram_cell[     341] = 32'h23871bb4;
    ram_cell[     342] = 32'h8c550e0f;
    ram_cell[     343] = 32'h8ac13b59;
    ram_cell[     344] = 32'hb6109a1b;
    ram_cell[     345] = 32'h80bb1e66;
    ram_cell[     346] = 32'h145a773c;
    ram_cell[     347] = 32'he8eb9a15;
    ram_cell[     348] = 32'hac631b41;
    ram_cell[     349] = 32'h84ef6c0a;
    ram_cell[     350] = 32'h1c7d3a9c;
    ram_cell[     351] = 32'h62b5b573;
    ram_cell[     352] = 32'h628b6ff4;
    ram_cell[     353] = 32'h6705c7b1;
    ram_cell[     354] = 32'ha1bdb151;
    ram_cell[     355] = 32'hcf40ef63;
    ram_cell[     356] = 32'h4eb51c01;
    ram_cell[     357] = 32'hab70fac7;
    ram_cell[     358] = 32'hbabcaec6;
    ram_cell[     359] = 32'hc7ae3652;
    ram_cell[     360] = 32'h64c81f38;
    ram_cell[     361] = 32'h846d0a87;
    ram_cell[     362] = 32'h4fb54152;
    ram_cell[     363] = 32'hf3e3a0c3;
    ram_cell[     364] = 32'hcd790ed1;
    ram_cell[     365] = 32'ha777dad5;
    ram_cell[     366] = 32'h7fa2183b;
    ram_cell[     367] = 32'h7c4da673;
    ram_cell[     368] = 32'hd97c83c1;
    ram_cell[     369] = 32'hc60bfd44;
    ram_cell[     370] = 32'h505402a7;
    ram_cell[     371] = 32'haf8d6023;
    ram_cell[     372] = 32'h523096b8;
    ram_cell[     373] = 32'h9befad0c;
    ram_cell[     374] = 32'hd30359e3;
    ram_cell[     375] = 32'h98ba90c0;
    ram_cell[     376] = 32'hc97a8ba4;
    ram_cell[     377] = 32'h2ebb1c49;
    ram_cell[     378] = 32'h9891ecf7;
    ram_cell[     379] = 32'h89973b86;
    ram_cell[     380] = 32'hf7e180ec;
    ram_cell[     381] = 32'hc4601887;
    ram_cell[     382] = 32'h563d36da;
    ram_cell[     383] = 32'h41b00c32;
    ram_cell[     384] = 32'ha4773e29;
    ram_cell[     385] = 32'hb265471c;
    ram_cell[     386] = 32'hb9218a97;
    ram_cell[     387] = 32'h2cf7f642;
    ram_cell[     388] = 32'hc4938215;
    ram_cell[     389] = 32'hbc141884;
    ram_cell[     390] = 32'hf60d0565;
    ram_cell[     391] = 32'h4ef78a24;
    ram_cell[     392] = 32'h4824bebc;
    ram_cell[     393] = 32'h9f2e6c40;
    ram_cell[     394] = 32'he0ad771f;
    ram_cell[     395] = 32'h66973958;
    ram_cell[     396] = 32'h7130611a;
    ram_cell[     397] = 32'hfffecbf6;
    ram_cell[     398] = 32'h618512e2;
    ram_cell[     399] = 32'hf92245ac;
    ram_cell[     400] = 32'h96974df1;
    ram_cell[     401] = 32'h94bd9337;
    ram_cell[     402] = 32'h56994807;
    ram_cell[     403] = 32'heb711500;
    ram_cell[     404] = 32'h36cf1544;
    ram_cell[     405] = 32'h6335ed1c;
    ram_cell[     406] = 32'h5fa03820;
    ram_cell[     407] = 32'hafbaa878;
    ram_cell[     408] = 32'h9f928387;
    ram_cell[     409] = 32'hf62daa2a;
    ram_cell[     410] = 32'hb35ef787;
    ram_cell[     411] = 32'hf8d39e36;
    ram_cell[     412] = 32'h898bc7cd;
    ram_cell[     413] = 32'hebe99110;
    ram_cell[     414] = 32'h2f137c5c;
    ram_cell[     415] = 32'h26c7018d;
    ram_cell[     416] = 32'h61ce28a5;
    ram_cell[     417] = 32'h0b4a2682;
    ram_cell[     418] = 32'hccb51607;
    ram_cell[     419] = 32'h95888111;
    ram_cell[     420] = 32'hf25ca604;
    ram_cell[     421] = 32'h12aa12ef;
    ram_cell[     422] = 32'h20f49505;
    ram_cell[     423] = 32'h0b58dd94;
    ram_cell[     424] = 32'hd6d56ddf;
    ram_cell[     425] = 32'hfe5460c3;
    ram_cell[     426] = 32'hf026023a;
    ram_cell[     427] = 32'h31212b11;
    ram_cell[     428] = 32'hbeb0d205;
    ram_cell[     429] = 32'h61d07aca;
    ram_cell[     430] = 32'he2a0c0a2;
    ram_cell[     431] = 32'h547e7e30;
    ram_cell[     432] = 32'h593b33c1;
    ram_cell[     433] = 32'h00636ad6;
    ram_cell[     434] = 32'h227a1223;
    ram_cell[     435] = 32'h1df2c16b;
    ram_cell[     436] = 32'h794c9906;
    ram_cell[     437] = 32'h77f918d3;
    ram_cell[     438] = 32'hd7e5319c;
    ram_cell[     439] = 32'h65f437d3;
    ram_cell[     440] = 32'had52f31e;
    ram_cell[     441] = 32'h9ed25a91;
    ram_cell[     442] = 32'hfef8e78f;
    ram_cell[     443] = 32'h9e08ecf2;
    ram_cell[     444] = 32'h818f0aba;
    ram_cell[     445] = 32'ha3a6a98f;
    ram_cell[     446] = 32'h04bddf0b;
    ram_cell[     447] = 32'h3d601a78;
    ram_cell[     448] = 32'h59a61093;
    ram_cell[     449] = 32'h04ab8a49;
    ram_cell[     450] = 32'h1b8937ec;
    ram_cell[     451] = 32'he6a40038;
    ram_cell[     452] = 32'h03fa8592;
    ram_cell[     453] = 32'he7a523d3;
    ram_cell[     454] = 32'hfd307558;
    ram_cell[     455] = 32'hdebcaa6a;
    ram_cell[     456] = 32'h9605160f;
    ram_cell[     457] = 32'h89ea2891;
    ram_cell[     458] = 32'hf64da302;
    ram_cell[     459] = 32'h76b3ed2f;
    ram_cell[     460] = 32'hee6fffdc;
    ram_cell[     461] = 32'hf5fa79a5;
    ram_cell[     462] = 32'h10470016;
    ram_cell[     463] = 32'hf5d22236;
    ram_cell[     464] = 32'ha43f8f0f;
    ram_cell[     465] = 32'hbc004f01;
    ram_cell[     466] = 32'hc96aaef0;
    ram_cell[     467] = 32'h514121d2;
    ram_cell[     468] = 32'h9d847ae8;
    ram_cell[     469] = 32'h0269768e;
    ram_cell[     470] = 32'hadba8737;
    ram_cell[     471] = 32'hd351c539;
    ram_cell[     472] = 32'h608e1cc8;
    ram_cell[     473] = 32'heb36fc06;
    ram_cell[     474] = 32'hd30f62bb;
    ram_cell[     475] = 32'h7266c1c2;
    ram_cell[     476] = 32'hcc475518;
    ram_cell[     477] = 32'hff04af83;
    ram_cell[     478] = 32'h2167e0ff;
    ram_cell[     479] = 32'h2bd5317c;
    ram_cell[     480] = 32'hf3a39fda;
    ram_cell[     481] = 32'hd02c5603;
    ram_cell[     482] = 32'h31b20e80;
    ram_cell[     483] = 32'h7282079b;
    ram_cell[     484] = 32'h05add105;
    ram_cell[     485] = 32'h1eeaa949;
    ram_cell[     486] = 32'h59a1ba1c;
    ram_cell[     487] = 32'h8400d987;
    ram_cell[     488] = 32'h2b57873f;
    ram_cell[     489] = 32'h2e714215;
    ram_cell[     490] = 32'hf52f0a23;
    ram_cell[     491] = 32'ha50c032d;
    ram_cell[     492] = 32'h941ab584;
    ram_cell[     493] = 32'h8e4f2ec6;
    ram_cell[     494] = 32'h455df895;
    ram_cell[     495] = 32'he2cbc402;
    ram_cell[     496] = 32'h0dda30a2;
    ram_cell[     497] = 32'h6eb8bb07;
    ram_cell[     498] = 32'h34b68fea;
    ram_cell[     499] = 32'h1697cfee;
    ram_cell[     500] = 32'hf1564ff0;
    ram_cell[     501] = 32'h92404a2f;
    ram_cell[     502] = 32'h582a5e82;
    ram_cell[     503] = 32'h6dfbd490;
    ram_cell[     504] = 32'h2d5566bf;
    ram_cell[     505] = 32'h846af710;
    ram_cell[     506] = 32'h7f8fc2e8;
    ram_cell[     507] = 32'hdb67d64e;
    ram_cell[     508] = 32'h961b6247;
    ram_cell[     509] = 32'hb4743d3c;
    ram_cell[     510] = 32'hcf79a7fd;
    ram_cell[     511] = 32'ha89c54d8;
    // src matrix B
    ram_cell[     512] = 32'hcd3a57e3;
    ram_cell[     513] = 32'hae39312e;
    ram_cell[     514] = 32'h2c691129;
    ram_cell[     515] = 32'h06bd3e43;
    ram_cell[     516] = 32'h23be9224;
    ram_cell[     517] = 32'hd4e3a778;
    ram_cell[     518] = 32'h76321322;
    ram_cell[     519] = 32'h688362c4;
    ram_cell[     520] = 32'h5e982c87;
    ram_cell[     521] = 32'ha7759da9;
    ram_cell[     522] = 32'hb0709ad4;
    ram_cell[     523] = 32'h8027987f;
    ram_cell[     524] = 32'h11addf09;
    ram_cell[     525] = 32'h9261244c;
    ram_cell[     526] = 32'h05353461;
    ram_cell[     527] = 32'h114bcb95;
    ram_cell[     528] = 32'h7bf4fcfe;
    ram_cell[     529] = 32'h35407dad;
    ram_cell[     530] = 32'hdc8675af;
    ram_cell[     531] = 32'hde2b6f57;
    ram_cell[     532] = 32'h467a546e;
    ram_cell[     533] = 32'ha8eca1d0;
    ram_cell[     534] = 32'h0d97628c;
    ram_cell[     535] = 32'h4c38438c;
    ram_cell[     536] = 32'h02239064;
    ram_cell[     537] = 32'hc40b7b06;
    ram_cell[     538] = 32'h87cfefa6;
    ram_cell[     539] = 32'he37197a0;
    ram_cell[     540] = 32'hae7a2621;
    ram_cell[     541] = 32'h7e995cfc;
    ram_cell[     542] = 32'h7a4a98ef;
    ram_cell[     543] = 32'h3ef881df;
    ram_cell[     544] = 32'hf1304336;
    ram_cell[     545] = 32'h737c22db;
    ram_cell[     546] = 32'h19ae0cf7;
    ram_cell[     547] = 32'h8b66d02d;
    ram_cell[     548] = 32'ha4352d17;
    ram_cell[     549] = 32'hc79f35d9;
    ram_cell[     550] = 32'h8dffd300;
    ram_cell[     551] = 32'h47b3cc71;
    ram_cell[     552] = 32'h3534250f;
    ram_cell[     553] = 32'h1461ec32;
    ram_cell[     554] = 32'h2ccfa14f;
    ram_cell[     555] = 32'h05bd2b86;
    ram_cell[     556] = 32'h3a9bf2ea;
    ram_cell[     557] = 32'h91d47366;
    ram_cell[     558] = 32'he000d0fc;
    ram_cell[     559] = 32'h8850674b;
    ram_cell[     560] = 32'hb1e06e7a;
    ram_cell[     561] = 32'h65c0c9c4;
    ram_cell[     562] = 32'hfb571e7e;
    ram_cell[     563] = 32'hc4517bbb;
    ram_cell[     564] = 32'h78b98121;
    ram_cell[     565] = 32'hf6e7e3fc;
    ram_cell[     566] = 32'hf1553cb6;
    ram_cell[     567] = 32'haf44a200;
    ram_cell[     568] = 32'h130c40fb;
    ram_cell[     569] = 32'he966109a;
    ram_cell[     570] = 32'hf4c13477;
    ram_cell[     571] = 32'h7532b6e8;
    ram_cell[     572] = 32'hd500282f;
    ram_cell[     573] = 32'hfcae77b5;
    ram_cell[     574] = 32'h0f799da3;
    ram_cell[     575] = 32'hc68b5e4d;
    ram_cell[     576] = 32'h5110f9fa;
    ram_cell[     577] = 32'hbf94f5ec;
    ram_cell[     578] = 32'h32b1f1e8;
    ram_cell[     579] = 32'h818d1b5d;
    ram_cell[     580] = 32'hec312908;
    ram_cell[     581] = 32'h0a1d382e;
    ram_cell[     582] = 32'h78df8919;
    ram_cell[     583] = 32'h59234837;
    ram_cell[     584] = 32'h011a4bdf;
    ram_cell[     585] = 32'h6961acae;
    ram_cell[     586] = 32'hb3ad4f3f;
    ram_cell[     587] = 32'h38e65234;
    ram_cell[     588] = 32'h0451268f;
    ram_cell[     589] = 32'h625117fc;
    ram_cell[     590] = 32'h74779060;
    ram_cell[     591] = 32'hf8d9938c;
    ram_cell[     592] = 32'hf5cd3901;
    ram_cell[     593] = 32'h923c7b72;
    ram_cell[     594] = 32'h12b3c034;
    ram_cell[     595] = 32'h80a8aa7f;
    ram_cell[     596] = 32'h516e716f;
    ram_cell[     597] = 32'hf359daa0;
    ram_cell[     598] = 32'h768ac36a;
    ram_cell[     599] = 32'h4f9976ea;
    ram_cell[     600] = 32'he41c8cad;
    ram_cell[     601] = 32'h97248d5a;
    ram_cell[     602] = 32'he570ed79;
    ram_cell[     603] = 32'hd5a837fa;
    ram_cell[     604] = 32'h9f89ad4b;
    ram_cell[     605] = 32'h15afc7de;
    ram_cell[     606] = 32'h304a6d20;
    ram_cell[     607] = 32'hcaa957dc;
    ram_cell[     608] = 32'he22e332e;
    ram_cell[     609] = 32'h82c4d280;
    ram_cell[     610] = 32'h97488fa1;
    ram_cell[     611] = 32'he94e2428;
    ram_cell[     612] = 32'h6fe4b3e4;
    ram_cell[     613] = 32'h96d85ed4;
    ram_cell[     614] = 32'h3d4d3829;
    ram_cell[     615] = 32'h0baa5a6f;
    ram_cell[     616] = 32'he3788eb0;
    ram_cell[     617] = 32'h871a3d5b;
    ram_cell[     618] = 32'he1fe0c01;
    ram_cell[     619] = 32'h4a7b7403;
    ram_cell[     620] = 32'h4afdd8c4;
    ram_cell[     621] = 32'hcf7cfedf;
    ram_cell[     622] = 32'h39da117b;
    ram_cell[     623] = 32'hd81a276a;
    ram_cell[     624] = 32'hd4006525;
    ram_cell[     625] = 32'h41717475;
    ram_cell[     626] = 32'h72a70e26;
    ram_cell[     627] = 32'hb41c6128;
    ram_cell[     628] = 32'h4e9f1c6c;
    ram_cell[     629] = 32'hba6485bd;
    ram_cell[     630] = 32'h4ab34f55;
    ram_cell[     631] = 32'h300ecab2;
    ram_cell[     632] = 32'hd16d1904;
    ram_cell[     633] = 32'hd71cd6e9;
    ram_cell[     634] = 32'he7c4e714;
    ram_cell[     635] = 32'he057c8c4;
    ram_cell[     636] = 32'h55be78c7;
    ram_cell[     637] = 32'h5a6f3516;
    ram_cell[     638] = 32'hd3bf41f5;
    ram_cell[     639] = 32'haf9d2be5;
    ram_cell[     640] = 32'h1a50eea1;
    ram_cell[     641] = 32'h265f5fd6;
    ram_cell[     642] = 32'h6ee2d8b0;
    ram_cell[     643] = 32'hc15b1e53;
    ram_cell[     644] = 32'hf4c80305;
    ram_cell[     645] = 32'h0c2a860f;
    ram_cell[     646] = 32'h58340f7b;
    ram_cell[     647] = 32'h0558390f;
    ram_cell[     648] = 32'h30a5f56d;
    ram_cell[     649] = 32'hfd91b839;
    ram_cell[     650] = 32'h47547c13;
    ram_cell[     651] = 32'hb26d3a2a;
    ram_cell[     652] = 32'h7d5f07f7;
    ram_cell[     653] = 32'hca3bc894;
    ram_cell[     654] = 32'hb238bfbe;
    ram_cell[     655] = 32'h1fd0ad50;
    ram_cell[     656] = 32'hf451e9d9;
    ram_cell[     657] = 32'h14b5167f;
    ram_cell[     658] = 32'h15865968;
    ram_cell[     659] = 32'hf27df7ac;
    ram_cell[     660] = 32'h2132a247;
    ram_cell[     661] = 32'hf2448fee;
    ram_cell[     662] = 32'h1a0e8414;
    ram_cell[     663] = 32'h94127148;
    ram_cell[     664] = 32'hd732a749;
    ram_cell[     665] = 32'h605cfa37;
    ram_cell[     666] = 32'h0801040d;
    ram_cell[     667] = 32'h9f23b01c;
    ram_cell[     668] = 32'h033f37ac;
    ram_cell[     669] = 32'h00e985c9;
    ram_cell[     670] = 32'h6b483b62;
    ram_cell[     671] = 32'h5bd7c299;
    ram_cell[     672] = 32'h2b756f82;
    ram_cell[     673] = 32'he20afe33;
    ram_cell[     674] = 32'h836be0c8;
    ram_cell[     675] = 32'hb7f8d7fb;
    ram_cell[     676] = 32'h9c8e2a8d;
    ram_cell[     677] = 32'h38cb0204;
    ram_cell[     678] = 32'h24a98754;
    ram_cell[     679] = 32'h024beeec;
    ram_cell[     680] = 32'heb25d211;
    ram_cell[     681] = 32'hdc0afc59;
    ram_cell[     682] = 32'hf1af61fc;
    ram_cell[     683] = 32'h0c9b7d68;
    ram_cell[     684] = 32'hd89efe98;
    ram_cell[     685] = 32'h15d0174b;
    ram_cell[     686] = 32'h9ec90789;
    ram_cell[     687] = 32'h0c87ceda;
    ram_cell[     688] = 32'h821c5470;
    ram_cell[     689] = 32'h6d520000;
    ram_cell[     690] = 32'h1d8fc639;
    ram_cell[     691] = 32'h28065c9d;
    ram_cell[     692] = 32'h72a2fd36;
    ram_cell[     693] = 32'h9b00298f;
    ram_cell[     694] = 32'h15d10897;
    ram_cell[     695] = 32'h6cb05ba3;
    ram_cell[     696] = 32'h6c9dfbd7;
    ram_cell[     697] = 32'h11f3d78f;
    ram_cell[     698] = 32'hf1d6e51a;
    ram_cell[     699] = 32'h42b8f590;
    ram_cell[     700] = 32'h15280459;
    ram_cell[     701] = 32'hec770cc1;
    ram_cell[     702] = 32'h44184227;
    ram_cell[     703] = 32'heb08e59c;
    ram_cell[     704] = 32'h3be9290b;
    ram_cell[     705] = 32'h28a56222;
    ram_cell[     706] = 32'hac35b671;
    ram_cell[     707] = 32'h08790b3f;
    ram_cell[     708] = 32'h55adb464;
    ram_cell[     709] = 32'hdf2f8ce5;
    ram_cell[     710] = 32'h1e6864bb;
    ram_cell[     711] = 32'hdfd933ca;
    ram_cell[     712] = 32'he6a59e88;
    ram_cell[     713] = 32'hfcab0197;
    ram_cell[     714] = 32'h0aeafa62;
    ram_cell[     715] = 32'h1fb2b443;
    ram_cell[     716] = 32'hcfdef149;
    ram_cell[     717] = 32'hc657e428;
    ram_cell[     718] = 32'hfda35dcb;
    ram_cell[     719] = 32'h9b35e61e;
    ram_cell[     720] = 32'h72b95f8b;
    ram_cell[     721] = 32'h0501c46e;
    ram_cell[     722] = 32'h013cc28e;
    ram_cell[     723] = 32'h3e810ef8;
    ram_cell[     724] = 32'hdc30ee72;
    ram_cell[     725] = 32'heac43659;
    ram_cell[     726] = 32'hdcf38f43;
    ram_cell[     727] = 32'he0aff351;
    ram_cell[     728] = 32'h0c1d9d1a;
    ram_cell[     729] = 32'hd95c8a83;
    ram_cell[     730] = 32'hfa862df0;
    ram_cell[     731] = 32'hf5048bba;
    ram_cell[     732] = 32'h7ac0c569;
    ram_cell[     733] = 32'h39a5a0af;
    ram_cell[     734] = 32'h8918d4b2;
    ram_cell[     735] = 32'h2be708c7;
    ram_cell[     736] = 32'h6971ec67;
    ram_cell[     737] = 32'h5c58b068;
    ram_cell[     738] = 32'h38ea2ce5;
    ram_cell[     739] = 32'h4cb7a999;
    ram_cell[     740] = 32'h9daba7e6;
    ram_cell[     741] = 32'hf46a330a;
    ram_cell[     742] = 32'hd9a81f19;
    ram_cell[     743] = 32'h53601ccc;
    ram_cell[     744] = 32'hd16d88a2;
    ram_cell[     745] = 32'hecb3d2fb;
    ram_cell[     746] = 32'h0c56da9a;
    ram_cell[     747] = 32'h9af68c3f;
    ram_cell[     748] = 32'hdd222e1e;
    ram_cell[     749] = 32'h8e1be0d7;
    ram_cell[     750] = 32'hcb10da72;
    ram_cell[     751] = 32'h4cc97a04;
    ram_cell[     752] = 32'h17a40453;
    ram_cell[     753] = 32'he0d9be3b;
    ram_cell[     754] = 32'hc6653998;
    ram_cell[     755] = 32'h63bd4b3f;
    ram_cell[     756] = 32'h1d992951;
    ram_cell[     757] = 32'hbffe5f0a;
    ram_cell[     758] = 32'h06633070;
    ram_cell[     759] = 32'h8c5eded1;
    ram_cell[     760] = 32'h2385aee6;
    ram_cell[     761] = 32'hd4b8969c;
    ram_cell[     762] = 32'hfa00b998;
    ram_cell[     763] = 32'h60abf34c;
    ram_cell[     764] = 32'heb439e70;
    ram_cell[     765] = 32'h2c52dd7a;
    ram_cell[     766] = 32'hf3125a81;
    ram_cell[     767] = 32'h6bf463f3;
end

endmodule

